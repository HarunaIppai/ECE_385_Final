module spawn_control(
	input  logic [2:0] 	Spawn0Data;
	input  logic [2:0] 	Spawn1Data;
	input  logic 		 	Spawn0State;
	input  logic 			Spawn1State;
	input  logic			SpawnReset;
	output logic [2:0]	Spawn_0;
	output logic [2:0]	Spawn_1;
);

	always_comb begin
			if(SpawnReset)
	end
endmodule 